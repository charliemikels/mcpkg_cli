module main

import mcpkg

fn main() {
	println('Hello World!')
}
